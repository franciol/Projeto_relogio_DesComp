LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;

ENTITY IO IS
    GENERIC (
        quantidadeBotao : NATURAL := 1
    );

    PORT (
        habilita : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
        RESET_IN : IN STD_LOGIC;
        saidaSW0,saidaSW1, RESET_OUT : OUT STD_LOGIC
    );
END ENTITY;

ARCHITECTURE FILSDELA OF IO IS
BEGIN
    saidaSW0 <= '1' WHEN (habilita(0) = '1') ELSE -- ATIVA SAIDA BASE DE TEMPO
    '0';
    
    saidaSW1 <= '1' WHEN (habilita(1) = '1') ELSE -- ATIVA SAIDA BASE DE TEMPO
    '0';

    RESET_OUT <= '1' WHEN (RESET_IN = '0') ELSE -- ATIVA RESET
    '0';
        
END ARCHITECTURE;